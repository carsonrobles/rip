package uart_pkg;

  parameter bit UART_START_BIT = 1'b0;
  parameter bit UART_STOP_BIT  = 1'b1;

endpackage
